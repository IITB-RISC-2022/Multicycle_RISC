library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_word is 
	port (s: in std_logic_vector(4 downto 0);
			ir: in std_logic_vector(15 downto 0);
			X: out std_logic_vector(35 downto 0));
end entity;

architecture Behave of control_word is
	type bits is array(0 to 27) of std_logic_vector(35 downto 0);
	signal control_bits : bits :=  (			"000000000000000000000000000000000000",
												"000101000000000000000110000000000001",
												"100000010000000000000000000010010000",
												"000000000000011000001000000011000000",
												"000000001001000000000000000000000000",
												"000000000000010000001000000011000000",
												"000000000000010010001000000011000000",
												"000000001111000000000000000000000000",
												"000000000000100000000000000011000000",
												"000001000000000000000000000000001000",
												"000000001110000000000000000000000000",
												"001010000000000000000000010000000000",
												"100000000000000000000000000000110000",
												"100001000000000000000000000000101010",
												"000000000110011010000000000011000000",
												"100000000000000000000000000000100010",
												"000000100000000000000000000000000100",
												"010010000000000000000000010100000000",
												"000000110000011000110000000010000000",
												"000000000000010000000011001000000000",
												"000000110000000000000000000000000100",
												"000000001110110110000011001000000000",
												"000000001110000000000010111000000000",
												"100000010000000000000000000010110000",
												"000000000000000000000000100000000000",
												"000000000000000000000000010000000000",
												"000000000000000000000001000000000000",
												"100000000000100000000000000000000000");
begin
	process(s, ir)
		variable temp_x : std_logic_vector(35 downto 0);
	begin
		temp_x := control_bits(to_integer(unsigned(s)));
		if s = "00011" then
			case ir(15 downto 12) is
				when "0010" =>
					temp_x(18 downto 15) := "1011";
				when others =>
					temp_x(18 downto 17) := "00";
			end case;
		end if;
		X <= temp_x;
	end process;
end architecture;