-- IITB-RISC-2022
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY control_word IS
	PORT (
		s : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		ir : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		X : OUT STD_LOGIC_VECTOR(33 DOWNTO 0));
END ENTITY;

ARCHITECTURE Behave OF control_word IS
	TYPE bits IS ARRAY(0 TO 28) OF STD_LOGIC_VECTOR(33 DOWNTO 0);
	SIGNAL control_bits : bits := (
	"0000000000000000000000000000000000",
	"0001010000000000000001100000000001",
	"1000000100000000000000000010010000",
	"0000000000000110000010000011000000",
	"0000000010010000000000000000000000",
	"0000000000000100000010000011000000",
	"0000000000000100100010000011000000",
	"0000000011110000000000000000000000",
	"0000000000001000000000000011000000",
	"0000010000000000000000000000001000",
	"0000000011100000000000000000000000",
	"0010100000000000000000000000000000",
	"1000000000000000000000000000110000",
	"1000010000000000000000000000101010",
	"0000000001100110100000000011000000",
	"1000000000000000000000000000100010",
	"0000001000000000000000000000000100",
	"0100100000000000000000000100000000",
	"0000001100000110001100000010000000",
	"0000000000000100000000110000000000",
	"0000001100000000000000000000000100",
	"0000000011101101100000110000000000",
	"0000000011100000000000101000000000",
	"1000000100000000000000000010110000",
	"0000000000000000000000001000000000",
	"0000000000000000000000000000000000",
	"0000000000000000000000010000000000",
	"1000000000001000000000000000000000",
	"0000000000010000000000000000000000");
BEGIN
	PROCESS (s, ir)
		VARIABLE temp_x : STD_LOGIC_VECTOR(33 DOWNTO 0);
	BEGIN
		temp_x := control_bits(to_integer(unsigned(s)));
		IF s = "00011" THEN
			CASE ir(15 DOWNTO 12) IS
				WHEN "0010" =>
					temp_x(16 DOWNTO 13) := "1011";
				WHEN OTHERS =>
					temp_x(16 DOWNTO 15) := "00";
			END CASE;
		END IF;

		IF s = "10011" OR s = "10101" THEN
			CASE ir(15 DOWNTO 12) IS
				WHEN "1000" =>
					temp_x(16 DOWNTO 13) := "1100";
				WHEN "1001" =>
					temp_x(16 DOWNTO 13) := "1100";
				WHEN OTHERS =>
					temp_x(16 DOWNTO 15) := "00";
			END CASE;
		END IF;
		X <= temp_x;
	END PROCESS;
END ARCHITECTURE;