library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_word is 
	port (s: in std_logic_vector(4 downto 0);
			ir: in std_logic_vector(15 downto 0);
			X: out std_logic_vector(34 downto 0));
end entity;

architecture Behave of control_word is
	type bits is array(0 to 26) of std_logic_vector(34 downto 0);
	signal control_bits : bits :=  ("00000000000000000000000000000000000",
												"00101000000000000000110000000000001",
											   "00000010000000000000000000010010000",
												"00000000000011000001000000011000000",
												"00000001001000000000000000000000000",
												"00000000000010000001000000011000000",
												"00000000000010010001000000011000000",
												"00000001111000000000000000000000000",
												"00000000000100000000000000011000000",
												"00001000000000000000000000000001000",
												"00000001110000000000000000000000000",
												"01010000000000000000000010000000000",
												"00000000000000000000000000000110000",
												"00001000000000000000000000000101010",
												"00000000110011010000000000011000000",
												"00000000000000000000000000000100010",
												"00000100000000000000000000000000100",
												"10010000000000000000000010100000000",
												"00000110000011000110000000010000000",
												"00000000000010100000011001000000000",
												"00000110000000000000000000000000100",
												"00000001110110110000011001000000000",
												"00000001110000000000010111000000000",
												"00000010000000000000000000010110000",
												"00000000000000000000000100000000000",
												"00000000000000000000000010000000000",
												"00000000000000000000001000000000000");
begin
	process(s, ir)
		variable temp_x : std_logic_vector(34 downto 0);
	begin
		temp_x := control_bits(to_integer(unsigned(s)));
		case ir(15 downto 12) is
			when "0001" =>
				temp_x(18 downto 17) := "00";
			when "0010" =>
				temp_x(18 downto 17) := "10";
			when others => 
				
		end case;
		X <= temp_x;
	end process;
end architecture;