-- IITB-RISC-2022
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_word is 
	port (s: in std_logic_vector(4 downto 0);
			ir: in std_logic_vector(15 downto 0);
			X: out std_logic_vector(33 downto 0));
end entity;

architecture Behave of control_word is
	type bits is array(0 to 27) of std_logic_vector(33 downto 0);
	signal control_bits : bits :=  (	"0000000000000000000000000000000000",
	"0001010000000000000001100000000001",
	"1000000100000000000000000010010000",
	"0000000000000110000010000011000000",
	"0000000010010000000000000000000000",
	"0000000000000100000010000011000000",
	"0000000000000100100010000011000000",
	"0000000011110000000000000000000000",
	"0000000000001000000000000011000000",
	"0000010000000000000000000000001000",
	"0000000011100000000000000000000000",
	"0010100000000000000000000000000000",
	"1000000000000000000000000000110000",
	"1000010000000000000000000000101010",
	"0000000001100110100000000011000000",
	"1000000000000000000000000000100010",
	"0000001000000000000000000000000100",
	"0100100000000000000000000100000000",
	"0000001100000110001100000010000000",
	"0000000000000100000000110000000000",
	"0000001100000000000000000000000100",
	"0000000011101101100000110000000000",
	"0000000011100000000000101000000000",
	"1000000100000000000000000010110000",
	"0000000000000000000000001000000000",
	"0000000000000000000000000000000000",
	"0000000000000000000000010000000000",
	"1000000000001000000000000000000000");
begin
	process(s, ir)
		variable temp_x : std_logic_vector(33 downto 0);
	begin
		temp_x := control_bits(to_integer(unsigned(s)));
		if s = "00011" then
			case ir(15 downto 12) is
				when "0010" =>
					temp_x(16 downto 13) := "1011";
				when others =>
					temp_x(16 downto 15) := "00";
			end case;
		end if;

		if s = "10011" or s = "10101" then
			case ir(15 downto 12) is
				when "1000" =>
					temp_x(16 downto 13) := "1100";
				when "1001" =>
					temp_x(16 downto 13) := "1100";
				when others =>
					temp_x(16 downto 15) := "00";
			end case;
		end if;
		X <= temp_x;
	end process;
end architecture;